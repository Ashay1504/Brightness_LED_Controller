LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY LED_BRIGHTNESS IS 
	PORT (
			LED_BR_EN : IN STD_LOGIC;
			IO_DATA   : INOUT std_logic_vector(15 downto 0)
			);
END LED_BRIGHTNESS;